//  This module is created by Mohamed Maged
//  Undergraduate ECE student, Alexandria university.


module BaudGen();

endmodule